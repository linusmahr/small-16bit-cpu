parameter SOMETHING = 16;

`define SOMETHING_2 3'h0